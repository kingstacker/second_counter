//************************************************
//  Filename      : second_counter.v                             
//  Author        : kingstacker                  
//  Company       : School                       
//  Email         : kingstacker_work@163.com     
//  Device        : Altera cyclone4 ep4ce6f17c8  
//  Description   : second_counter;key0:stop and begin;
//                  key1:recording;
//                  key2:order print;                             
//************************************************
module  second_counter_top (
/*i*/   input    wire    clk              ,
        input    wire    rst_n            ,
        input    wire    key0             , //stop&begin;
        input    wire    key1             , //recording key;
        input    wire    key2             , //order print;
/*o*/   output   wire                  ,
        output   wire     
);




endmodule