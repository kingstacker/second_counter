//************************************************
//  Filename      : sco.v                             
//  Author        : kingstacker                  
//  Company       : School                       
//  Email         : kingstacker_work@163.com     
//  Device        : Altera cyclone4 ep4ce6f17c8  
//  Description   :                              
//************************************************
module  sco (
/*i*/   input    wire              clk                 ,
        input    wire              rst_n               ,
        input    wire              key_bs              , //begin and stop;
        input    wire              key_rec             , //recording;
        input    wire              key_dis             , //display the value;
/*o*/   output   wire    [47:0]    dout        
);




endmodule